module and_gate(
  input bit [3:0] a,b,
  output bit [3:0] y
);
  
  assign y = a & b;
  
  
endmodule